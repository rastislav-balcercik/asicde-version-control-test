entity new_entity_vhd is

-- new comment

end entity new_entity_vhd;


testchange