entity new_entity_vhd is

end entity new_entity_vhd;