entity testentity1_vhd is

end entity testentity1_vhd;