entity asd_vhd is

end entity asd_vhd;