entity entity1_vhd is

end entity entity1_vhd;